module mem
(
    input wire x,
    output wire nx
);
assign x = ~nx;
endmodule
